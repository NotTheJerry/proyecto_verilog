module Compuerta_AND ( input a, input b, output salida );

	assign salida = a & b;

endmodule
